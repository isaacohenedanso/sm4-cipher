LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor_four IS
	PORT (
		INPT_A, INPT_B, INPT_C, INPT_D : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END xor_four;

ARCHITECTURE Behavioral OF xor_four IS

BEGIN
	OUTP <= INPT_A XOR INPT_B XOR INPT_C XOR INPT_D;
END Behavioral;