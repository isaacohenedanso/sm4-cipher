LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux1 IS
	PORT (
		SEL : IN STD_LOGIC;
		INPT_A, INPT_B : IN STD_LOGIC;
		OUTP : OUT STD_LOGIC
	);
END mux1;

ARCHITECTURE Behavioral OF mux1 IS

BEGIN
	WITH SEL SELECT
		OUTP <= INPT_A WHEN '0',
		INPT_B WHEN '1',
		'Z' WHEN OTHERS;
END Behavioral;