LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux32 IS
	PORT (
		SEL : IN STD_LOGIC;
		INPT_A, INPT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END mux32;

ARCHITECTURE Behavioral OF mux32 IS

BEGIN
	WITH SEL SELECT
		OUTP <= INPT_A WHEN '0',
		INPT_B WHEN '1',
		(OTHERS => '0') WHEN OTHERS;
END Behavioral;