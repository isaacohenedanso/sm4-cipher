LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor_three IS
	PORT (
		INPT_A, INPT_B, INPT_C : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END xor_three;

ARCHITECTURE Behavioral OF xor_three IS

BEGIN
	OUTP <= INPT_A XOR INPT_B XOR INPT_C;
END Behavioral;