LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY regi IS
	PORT (
		CLK, LOAD, RST : IN STD_LOGIC;
		D : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		Q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END regi;

ARCHITECTURE Behavioral OF regi IS
BEGIN
	PROCESS (CLK, RST) IS
	BEGIN
		IF (RST = '1') THEN
			Q <= "000000";
		ELSIF (rising_edge(CLK)) THEN
			IF (LOAD = '1') THEN
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;