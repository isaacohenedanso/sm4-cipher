LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Datapath IS
	PORT (
		INPUTTEXT, MASTERKEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		OUTPUTTEXT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		ENC_DEC, CLK, CLR, MKLOAD, ILOAD, XLOAD, MUXSEL1, MUXSEL2, MUXSEL3, MUXSEL4, WRITE_EN, OUTEN : IN STD_LOGIC;
		ILT32 : OUT STD_LOGIC
	);
END Datapath;

ARCHITECTURE Behavioral OF Datapath IS
	COMPONENT CounterAndRam IS
		PORT (
			WRITE_EN, ENC_DEC, CLK, RST, ILOAD, MUXSEL4 : IN STD_LOGIC;
			ILT32 : OUT STD_LOGIC;
			ROUNDKEY_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			ROUNDKEY_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			COUNT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT EncryptionDecryptionUnit IS
		PORT (
			XLOAD, CLK, MUXSEL3, OUTEN : IN STD_LOGIC;
			INPUTTEXT : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			ROUNDKEY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTPUTTEXT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT KeyExpansionUnit IS
		PORT (
			MKLOAD, CLK, MUXSEL1, MUXSEL2 : IN STD_LOGIC;
			MASTERKEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			ROUNDKEY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL ADDRESS_OF_ROM : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL GENERATED_ROUND_KEYS, KEYS_FROM_RAM : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	KeyExpansionUnit0 : KeyExpansionUnit PORT MAP(
		MKLOAD => MKLOAD,
		CLK => CLK,
		MASTERKEY => MASTERKEY,
		ADDRESS => ADDRESS_OF_ROM,
		MUXSEL1 => MUXSEL1,
		MUXSEL2 => MUXSEL2,
		ROUNDKEY => GENERATED_ROUND_KEYS
	);
	EncryptionDecryptionUnit0 : EncryptionDecryptionUnit PORT MAP(
		XLOAD => XLOAD,
		CLK => CLK,
		MUXSEL3 => MUXSEL3,
		OUTEN => OUTEN,
		INPUTTEXT => INPUTTEXT,
		ROUNDKEY => KEYS_FROM_RAM,
		OUTPUTTEXT => OUTPUTTEXT
	);
	CounterAndRam0 : CounterAndRam PORT MAP(
		WRITE_EN => WRITE_EN,
		ENC_DEC => ENC_DEC,
		CLK => CLK,
		RST => CLR,
		ILOAD => ILOAD,
		MUXSEL4 => MUXSEL4,
		ILT32 => ILT32,
		ROUNDKEY_IN => GENERATED_ROUND_KEYS,
		ROUNDKEY_OUT => KEYS_FROM_RAM,
		COUNT => ADDRESS_OF_ROM
	);

END Behavioral;