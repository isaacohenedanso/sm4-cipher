LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY KeyExpansionUnit IS
	PORT (
		MKLOAD, CLK, MUXSEL1, MUXSEL2 : IN STD_LOGIC;
		MASTERKEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		ROUNDKEY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END KeyExpansionUnit;

ARCHITECTURE Behavioral OF KeyExpansionUnit IS
	COMPONENT mux128 IS
		PORT (
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			SEL : IN STD_LOGIC;
			OUTP : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT reg128 IS
		PORT (
			CLK, LOAD : IN STD_LOGIC;
			D : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			Q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_four IS
		PORT (
			INPT_A, INPT_B, INPT_C, INPT_D : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_two IS
		PORT (
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT rom IS
		PORT (
			INPT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT sbox IS
		PORT (
			INPT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT mux96 IS
		PORT (
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(95 DOWNTO 0);
			SEL : IN STD_LOGIC;
			OUTP : OUT STD_LOGIC_VECTOR(95 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT mux32 IS
		PORT (
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			SEL : IN STD_LOGIC;
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_three IS
		PORT (
			INPT_A, INPT_B, INPT_C : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL FROMREGMK, FROMMUX128, NEXTINPT : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL FROMMUX96, K : STD_LOGIC_VECTOR(95 DOWNTO 0);
	SIGNAL FROMSBOXES, FROMXOR2_0, TOSBOXES, CIRC_SHIFT13, CIRC_SHIFT23, FROMROM, FROMXOR4_0, FROMXOR4_1, K0, K1, K2, K3, FROMMUX32_1, FROMXOR3_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL FROMSBOX0, FROMSBOX1, FROMSBOX2, FROMSBOX3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
	FROMSBOXES <= FROMSBOX0 & FROMSBOX1 & FROMSBOX2 & FROMSBOX3;
	CIRC_SHIFT13 <= FROMSBOXES(18 DOWNTO 0) & FROMSBOXES(31 DOWNTO 19);
	CIRC_SHIFT23 <= FROMSBOXES(8 DOWNTO 0) & FROMSBOXES(31 DOWNTO 9);
	k <= K1 & K2 & K3;
	NEXTINPT <= FROMMUX96(95 DOWNTO 0) & FROMXOR2_0;
	ROUNDKEY <= FROMXOR2_0;
	mux0 : mux128 PORT MAP(
		INPT_A => MASTERKEY,
		INPT_B => NEXTINPT,
		SEL => MUXSEL1,
		OUTP => FROMMUX128
	);
	regMK : reg128 PORT MAP(
		CLK => CLK,
		LOAD => MKLOAD,
		D => FROMMUX128,
		Q => FROMREGMK
	);
	romCK : rom PORT MAP(
		INPT => ADDRESS,
		OUTP => FROMROM
	);
	xor4_0 : xor_four PORT MAP(
		INPT_A => FROMREGMK(95 DOWNTO 64),
		INPT_B => FROMREGMK(63 DOWNTO 32),
		INPT_C => FROMREGMK(31 DOWNTO 0),
		INPT_D => FROMROM,
		OUTP => FROMXOR4_0
	);
	xor2_0 : xor_two PORT MAP(
		INPT_A => x"A3B1BAC6",
		INPT_B => FROMREGMK(127 DOWNTO 96),
		OUTP => K0
	);
	xor2_1 : xor_two PORT MAP(
		INPT_A => x"56AA3350",
		INPT_B => FROMREGMK(95 DOWNTO 64),
		OUTP => K1
	);
	xor2_2 : xor_two PORT MAP(
		INPT_A => x"677D9197",
		INPT_B => FROMREGMK(63 DOWNTO 32),
		OUTP => K2
	);
	xor2_3 : xor_two PORT MAP(
		INPT_A => x"B27022DC",
		INPT_B => FROMREGMK(31 DOWNTO 0),
		OUTP => K3
	);
	muxtosbox : mux32 PORT MAP(
		INPT_A => FROMXOR4_0,
		INPT_B => FROMXOR4_1,
		SEL => MUXSEL2,
		OUTP => TOSBOXES
	);
	xor4_1 : xor_four PORT MAP(
		INPT_A => K1,
		INPT_B => K2,
		INPT_C => K3,
		INPT_D => FROMROM,
		OUTP => FROMXOR4_1
	);
	sbox0 : sbox PORT MAP(
		INPT => TOSBOXES(31 DOWNTO 24),
		OUTP => FROMSBOX0
	);
	sbox1 : sbox PORT MAP(
		INPT => TOSBOXES(23 DOWNTO 16),
		OUTP => FROMSBOX1
	);
	sbox2 : sbox PORT MAP(
		INPT => TOSBOXES(15 DOWNTO 8),
		OUTP => FROMSBOX2
	);
	sbox3 : sbox PORT MAP(
		INPT => TOSBOXES(7 DOWNTO 0),
		OUTP => FROMSBOX3
	);
	mux32_1 : MUX32 PORT MAP(
		INPT_A => FROMREGMK(127 DOWNTO 96),
		INPT_B => K0,
		SEL => MUXSEL2,
		OUTP => FROMMUX32_1
	);
	mux96_0 : mux96 PORT MAP(
		INPT_A => FROMREGMK(95 DOWNTO 0),
		INPT_B => K,
		SEL => MUXSEL2,
		OUTP => FROMMUX96
	);
	xor3_0 : xor_three PORT MAP(
		INPT_A => FROMSBOXES,
		INPT_B => CIRC_SHIFT13,
		INPT_C => CIRC_SHIFT23,
		OUTP => FROMXOR3_0
	);
	xor2_5 : xor_two PORT MAP(
		INPT_A => FROMXOR3_0,
		INPT_B => FROMMUX32_1,
		OUTP => FROMXOR2_0
	);

END Behavioral;