LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux3 IS
	PORT (
		SEL : IN STD_LOGIC;
		INPT_A, INPT_B : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END mux3;

ARCHITECTURE Behavioral OF mux3 IS

BEGIN
	WITH SEL SELECT
		OUTP <= INPT_A WHEN '0',
		INPT_B WHEN '1',
		"ZZZ" WHEN OTHERS;
END Behavioral;