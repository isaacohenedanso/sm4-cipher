LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux128 IS
	PORT (
		SEL : IN STD_LOGIC;
		INPT_A, INPT_B : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END mux128;

ARCHITECTURE Behavioral OF mux128 IS

BEGIN
	WITH SEL SELECT
		OUTP <= INPT_A WHEN '0',
		INPT_B WHEN '1',
		(OTHERS => '0') WHEN OTHERS;
END Behavioral;