LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--
ENTITY adder IS
	PORT (
		INPT : IN unsigned(5 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END adder;

ARCHITECTURE Behavioral OF adder IS
BEGIN
	OUTP <= STD_LOGIC_VECTOR(INPT + 1);
END Behavioral;