LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux96 IS
	PORT (
		SEL : IN STD_LOGIC;
		INPT_A, INPT_B : IN STD_LOGIC_VECTOR(95 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(95 DOWNTO 0)
	);
END mux96;

ARCHITECTURE Behavioral OF mux96 IS

BEGIN
	WITH SEL SELECT
		OUTP <= INPT_A WHEN '0',
		INPT_B WHEN '1',
		(OTHERS => '0') WHEN OTHERS;
END Behavioral;