library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sbox is
	port(
		INPT: in std_logic_vector(7 downto 0);
		OUTP: out std_logic_vector(7 downto 0)
	);
end sbox;

architecture Behavioral of sbox is

begin
	with INPT select 
		OUTP <= x"D6" when x"00",
				x"90" when x"01",
				x"E9" when x"02",
				x"FE" when x"03",
				x"CC" when x"04",
				x"E1" when x"05",
				x"3D" when x"06",
				x"B7" when x"07",
				x"16" when x"08",
				x"B6" when x"09",
				x"14" when x"0A",
				x"C2" when x"0B",
				x"28" when x"0C",
				x"FB" when x"0D",
				x"2C" when x"0E",
				x"05" when x"0F",
				x"2B" when x"10",
				x"67" when x"11",
				x"9A" when x"12",
				x"76" when x"13",
				x"2A" when x"14",
				x"BE" when x"15",
				x"04" when x"16",
				x"C3" when x"17",
				x"AA" when x"18",
				x"44" when x"19",
				x"13" when x"1A",
				x"26" when x"1B",
				x"49" when x"1C",
				x"86" when x"1D",
				x"06" when x"1E",
				x"99" when x"1F",
				x"9C" when x"20",
				x"42" when x"21",
				x"50" when x"22",
				x"F4" when x"23",
				x"91" when x"24",
				x"EF" when x"25",
				x"98" when x"26",
				x"71" when x"27",
				x"33" when x"28",
				x"54" when x"29",
				x"0B" when x"2A",
				x"43" when x"2B",
				x"ED" when x"2C",
				x"CF" when x"2D",
				x"AC" when x"2E",
				x"62" when x"2F",
				x"E4" when x"30",
				x"B3" when x"31",
				x"1C" when x"32",
				x"A9" when x"33",
				x"C9" when x"34",
				x"08" when x"35",
				x"E8" when x"36",
				x"95" when x"37",
				x"80" when x"38",
				x"DF" when x"39",
				x"94" when x"3A",
				x"FA" when x"3B",
				x"75" when x"3C",
				x"8F" when x"3D",
				x"3F" when x"3E",
				x"A6" when x"3F",
				x"47" when x"40",
				x"07" when x"41",
				x"A7" when x"42",
				x"FC" when x"43",
				x"F3" when x"44",
				x"73" when x"45",
				x"17" when x"46",
				x"BA" when x"47",
				x"83" when x"48",
				x"59" when x"49",
				x"3C" when x"4A",
				x"19" when x"4B",
				x"E6" when x"4C",
				x"85" when x"4D",
				x"4F" when x"4E",
				x"A8" when x"4F",
				x"68" when x"50",
				x"6B" when x"51",
				x"81" when x"52",
				x"B2" when x"53",
				x"71" when x"54",
				x"64" when x"55",
				x"DA" when x"56",
				x"8B" when x"57",
				x"F8" when x"58",
				x"EB" when x"59",
				x"0F" when x"5A",
				x"4B" when x"5B",
				x"70" when x"5C",
				x"56" when x"5D",
				x"9D" when x"5E",
				x"35" when x"5F",
				x"1E" when x"60",
				x"24" when x"61",
				x"0E" when x"62",
				x"5E" when x"63",
				x"63" when x"64",
				x"58" when x"65",
				x"D1" when x"66",
				x"A2" when x"67",
				x"25" when x"68",
				x"22" when x"69",
				x"7C" when x"6A",
				x"3B" when x"6B",
				x"01" when x"6C",
				x"21" when x"6D",
				x"78" when x"6E",
				x"87" when x"6F",
				x"D4" when x"70",
				x"00" when x"71",
				x"46" when x"72",
				x"57" when x"73",
				x"9F" when x"74",
				x"D3" when x"75",
				x"27" when x"76",
				x"52" when x"77",
				x"4C" when x"78",
				x"36" when x"79",
				x"02" when x"7A",
				x"E7" when x"7B",
				x"A0" when x"7C",
				x"C4" when x"7D",
				x"C8" when x"7E",
				x"9E" when x"7F",
				x"EA" when x"80",
				x"B1" when x"81",
				x"8A" when x"82",
				x"D2" when x"83",
				x"40" when x"84",
				x"C7" when x"85",
				x"38" when x"86",
				x"B5" when x"87",
				x"A3" when x"88",
				x"F7" when x"89",
				x"F2" when x"8A",
				x"CE" when x"8B",
				x"F9" when x"8C",
				x"61" when x"8D",
				x"15" when x"8E",
				x"A1" when x"8F",
				x"E0" when x"90",
				x"AE" when x"91",
				x"5D" when x"92",
				x"A4" when x"93",
				x"9B" when x"94",
				x"34" when x"95",
				x"1A" when x"96",
				x"55" when x"97",
				x"AD" when x"98",
				x"93" when x"99",
				x"32" when x"9A",
				x"30" when x"9B",
				x"F5" when x"9C",
				x"8C" when x"9D",
				x"B1" when x"9E",
				x"E3" when x"9F",
				x"1D" when x"A0",
				x"F6" when x"A1",
				x"E2" when x"A2",
				x"2E" when x"A3",
				x"82" when x"A4",
				x"66" when x"A5",
				x"CA" when x"A6",
				x"60" when x"A7",
				x"C0" when x"A8",
				x"29" when x"A9",
				x"23" when x"AA",
				x"AB" when x"AB",
				x"0D" when x"AC",
				x"53" when x"AD",
				x"4E" when x"AE",
				x"6F" when x"AF",
				x"D5" when x"B0",
				x"DB" when x"B1",
				x"37" when x"B2",
				x"45" when x"B3",
				x"DE" when x"B4",
				x"FD" when x"B5",
				x"8E" when x"B6",
				x"2F" when x"B7",
				x"03" when x"B8",
				x"FF" when x"B9",
				x"6A" when x"BA",
				x"72" when x"BB",
				x"6D" when x"BC",
				x"6C" when x"BD",
				x"5B" when x"BE",
				x"51" when x"BF",
				x"8D" when x"C0",
				x"1B" when x"C1",
				x"AF" when x"C2",
				x"92" when x"C3",
				x"BB" when x"C4",
				x"DD" when x"C5",
				x"BC" when x"C6",
				x"7F" when x"C7",
				x"11" when x"C8",
				x"D9" when x"C9",
				x"5C" when x"CA",
				x"41" when x"CB",
				x"1F" when x"CC",
				x"10" when x"CD",
				x"5A" when x"CE",
				x"D8" when x"CF",
				x"0A" when x"D0",
				x"C1" when x"D1",
				x"31" when x"D2",
				x"88" when x"D3",
				x"A5" when x"D4",
				x"CD" when x"D5",
				x"7B" when x"D6",
				x"BD" when x"D7",
				x"2D" when x"D8",
				x"74" when x"D9",
				x"D0" when x"DA",
				x"12" when x"DB",
				x"B8" when x"DC",
				x"E5" when x"DD",
				x"B4" when x"DE",
				x"B0" when x"DF",
				x"89" when x"E0",
				x"69" when x"E1",
				x"97" when x"E2",
				x"4A" when x"E3",
				x"0C" when x"E4",
				x"96" when x"E5",
				x"77" when x"E6",
				x"7E" when x"E7",
				x"65" when x"E8",
				x"B9" when x"E9",
				x"F1" when x"EA",
				x"09" when x"EB",
				x"C5" when x"EC",
				x"6E" when x"ED",
				x"C6" when x"EE",
				x"84" when x"EF",
				x"18" when x"F0",
				x"F0" when x"F1",
				x"7D" when x"F2",
				x"EC" when x"F3",
				x"3A" when x"F4",
				x"DC" when x"F5",
				x"4D" when x"F6",
				x"20" when x"F7",
				x"79" when x"F8",
				x"EE" when x"F9",
				x"5F" when x"FA",
				x"3E" when x"FB",
				x"D7" when x"FC",
				x"CB" when x"FD",
				x"39" when x"FE",
				x"48" when x"FF",
				(others => '0') when others;
	
end Behavioral;

