LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY reg128 IS
	PORT (
		CLK, LOAD : IN STD_LOGIC;
		D : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		Q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END reg128;

ARCHITECTURE Behavioral OF reg128 IS
BEGIN
	PROCESS (CLK) IS
	BEGIN
		IF (rising_edge(CLK)) THEN
			IF (LOAD = '1') THEN
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;