LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor_two IS
	PORT (
		INPT_A, INPT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END xor_two;

ARCHITECTURE Behavioral OF xor_two IS

BEGIN
	OUTP <= INPT_A XOR INPT_B;
END Behavioral;