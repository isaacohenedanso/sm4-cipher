LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY xor2 IS
	PORT (
		INPT_A, INPT_B : IN STD_LOGIC_VEC
		TOR(31 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END xor2;

ARCHITECTURE Behavioral OF xor2 IS

BEGIN
	OUTP <= INPT_A XOR INPT_B;
END Behavioral;