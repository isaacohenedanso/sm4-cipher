LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--
ENTITY substractor IS
	PORT (
		INPT : IN unsigned(4 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END substractor;

ARCHITECTURE Behavioral OF substractor IS
BEGIN
	OUTP <= STD_LOGIC_VECTOR(31 - INPT);
END Behavioral;