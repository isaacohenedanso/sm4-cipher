LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY sbox IS
	PORT (
		INPT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END sbox;

ARCHITECTURE Behavioral OF sbox IS

BEGIN
	WITH INPT SELECT
		OUTP <= x"D6" WHEN x"00",
		x"90" WHEN x"01",
		x"E9" WHEN x"02",
		x"FE" WHEN x"03",
		x"CC" WHEN x"04",
		x"E1" WHEN x"05",
		x"3D" WHEN x"06",
		x"B7" WHEN x"07",
		x"16" WHEN x"08",
		x"B6" WHEN x"09",
		x"14" WHEN x"0A",
		x"C2" WHEN x"0B",
		x"28" WHEN x"0C",
		x"FB" WHEN x"0D",
		x"2C" WHEN x"0E",
		x"05" WHEN x"0F",
		x"2B" WHEN x"10",
		x"67" WHEN x"11",
		x"9A" WHEN x"12",
		x"76" WHEN x"13",
		x"2A" WHEN x"14",
		x"BE" WHEN x"15",
		x"04" WHEN x"16",
		x"C3" WHEN x"17",
		x"AA" WHEN x"18",
		x"44" WHEN x"19",
		x"13" WHEN x"1A",
		x"26" WHEN x"1B",
		x"49" WHEN x"1C",
		x"86" WHEN x"1D",
		x"06" WHEN x"1E",
		x"99" WHEN x"1F",
		x"9C" WHEN x"20",
		x"42" WHEN x"21",
		x"50" WHEN x"22",
		x"F4" WHEN x"23",
		x"91" WHEN x"24",
		x"EF" WHEN x"25",
		x"98" WHEN x"26",
		x"7A" WHEN x"27",
		x"33" WHEN x"28",
		x"54" WHEN x"29",
		x"0B" WHEN x"2A",
		x"43" WHEN x"2B",
		x"ED" WHEN x"2C",
		x"CF" WHEN x"2D",
		x"AC" WHEN x"2E",
		x"62" WHEN x"2F",
		x"E4" WHEN x"30",
		x"B3" WHEN x"31",
		x"1C" WHEN x"32",
		x"A9" WHEN x"33",
		x"C9" WHEN x"34",
		x"08" WHEN x"35",
		x"E8" WHEN x"36",
		x"95" WHEN x"37",
		x"80" WHEN x"38",
		x"DF" WHEN x"39",
		x"94" WHEN x"3A",
		x"FA" WHEN x"3B",
		x"75" WHEN x"3C",
		x"8F" WHEN x"3D",
		x"3F" WHEN x"3E",
		x"A6" WHEN x"3F",
		x"47" WHEN x"40",
		x"07" WHEN x"41",
		x"A7" WHEN x"42",
		x"FC" WHEN x"43",
		x"F3" WHEN x"44",
		x"73" WHEN x"45",
		x"17" WHEN x"46",
		x"BA" WHEN x"47",
		x"83" WHEN x"48",
		x"59" WHEN x"49",
		x"3C" WHEN x"4A",
		x"19" WHEN x"4B",
		x"E6" WHEN x"4C",
		x"85" WHEN x"4D",
		x"4F" WHEN x"4E",
		x"A8" WHEN x"4F",
		x"68" WHEN x"50",
		x"6B" WHEN x"51",
		x"81" WHEN x"52",
		x"B2" WHEN x"53",
		x"71" WHEN x"54",
		x"64" WHEN x"55",
		x"DA" WHEN x"56",
		x"8B" WHEN x"57",
		x"F8" WHEN x"58",
		x"EB" WHEN x"59",
		x"0F" WHEN x"5A",
		x"4B" WHEN x"5B",
		x"70" WHEN x"5C",
		x"56" WHEN x"5D",
		x"9D" WHEN x"5E",
		x"35" WHEN x"5F",
		x"1E" WHEN x"60",
		x"24" WHEN x"61",
		x"0E" WHEN x"62",
		x"5E" WHEN x"63",
		x"63" WHEN x"64",
		x"58" WHEN x"65",
		x"D1" WHEN x"66",
		x"A2" WHEN x"67",
		x"25" WHEN x"68",
		x"22" WHEN x"69",
		x"7C" WHEN x"6A",
		x"3B" WHEN x"6B",
		x"01" WHEN x"6C",
		x"21" WHEN x"6D",
		x"78" WHEN x"6E",
		x"87" WHEN x"6F",
		x"D4" WHEN x"70",
		x"00" WHEN x"71",
		x"46" WHEN x"72",
		x"57" WHEN x"73",
		x"9F" WHEN x"74",
		x"D3" WHEN x"75",
		x"27" WHEN x"76",
		x"52" WHEN x"77",
		x"4C" WHEN x"78",
		x"36" WHEN x"79",
		x"02" WHEN x"7A",
		x"E7" WHEN x"7B",
		x"A0" WHEN x"7C",
		x"C4" WHEN x"7D",
		x"C8" WHEN x"7E",
		x"9E" WHEN x"7F",
		x"EA" WHEN x"80",
		x"BF" WHEN x"81",
		x"8A" WHEN x"82",
		x"D2" WHEN x"83",
		x"40" WHEN x"84",
		x"C7" WHEN x"85",
		x"38" WHEN x"86",
		x"B5" WHEN x"87",
		x"A3" WHEN x"88",
		x"F7" WHEN x"89",
		x"F2" WHEN x"8A",
		x"CE" WHEN x"8B",
		x"F9" WHEN x"8C",
		x"61" WHEN x"8D",
		x"15" WHEN x"8E",
		x"A1" WHEN x"8F",
		x"E0" WHEN x"90",
		x"AE" WHEN x"91",
		x"5D" WHEN x"92",
		x"A4" WHEN x"93",
		x"9B" WHEN x"94",
		x"34" WHEN x"95",
		x"1A" WHEN x"96",
		x"55" WHEN x"97",
		x"AD" WHEN x"98",
		x"93" WHEN x"99",
		x"32" WHEN x"9A",
		x"30" WHEN x"9B",
		x"F5" WHEN x"9C",
		x"8C" WHEN x"9D",
		x"B1" WHEN x"9E",
		x"E3" WHEN x"9F",
		x"1D" WHEN x"A0",
		x"F6" WHEN x"A1",
		x"E2" WHEN x"A2",
		x"2E" WHEN x"A3",
		x"82" WHEN x"A4",
		x"66" WHEN x"A5",
		x"CA" WHEN x"A6",
		x"60" WHEN x"A7",
		x"C0" WHEN x"A8",
		x"29" WHEN x"A9",
		x"23" WHEN x"AA",
		x"AB" WHEN x"AB",
		x"0D" WHEN x"AC",
		x"53" WHEN x"AD",
		x"4E" WHEN x"AE",
		x"6F" WHEN x"AF",
		x"D5" WHEN x"B0",
		x"DB" WHEN x"B1",
		x"37" WHEN x"B2",
		x"45" WHEN x"B3",
		x"DE" WHEN x"B4",
		x"FD" WHEN x"B5",
		x"8E" WHEN x"B6",
		x"2F" WHEN x"B7",
		x"03" WHEN x"B8",
		x"FF" WHEN x"B9",
		x"6A" WHEN x"BA",
		x"72" WHEN x"BB",
		x"6D" WHEN x"BC",
		x"6C" WHEN x"BD",
		x"5B" WHEN x"BE",
		x"51" WHEN x"BF",
		x"8D" WHEN x"C0",
		x"1B" WHEN x"C1",
		x"AF" WHEN x"C2",
		x"92" WHEN x"C3",
		x"BB" WHEN x"C4",
		x"DD" WHEN x"C5",
		x"BC" WHEN x"C6",
		x"7F" WHEN x"C7",
		x"11" WHEN x"C8",
		x"D9" WHEN x"C9",
		x"5C" WHEN x"CA",
		x"41" WHEN x"CB",
		x"1F" WHEN x"CC",
		x"10" WHEN x"CD",
		x"5A" WHEN x"CE",
		x"D8" WHEN x"CF",
		x"0A" WHEN x"D0",
		x"C1" WHEN x"D1",
		x"31" WHEN x"D2",
		x"88" WHEN x"D3",
		x"A5" WHEN x"D4",
		x"CD" WHEN x"D5",
		x"7B" WHEN x"D6",
		x"BD" WHEN x"D7",
		x"2D" WHEN x"D8",
		x"74" WHEN x"D9",
		x"D0" WHEN x"DA",
		x"12" WHEN x"DB",
		x"B8" WHEN x"DC",
		x"E5" WHEN x"DD",
		x"B4" WHEN x"DE",
		x"B0" WHEN x"DF",
		x"89" WHEN x"E0",
		x"69" WHEN x"E1",
		x"97" WHEN x"E2",
		x"4A" WHEN x"E3",
		x"0C" WHEN x"E4",
		x"96" WHEN x"E5",
		x"77" WHEN x"E6",
		x"7E" WHEN x"E7",
		x"65" WHEN x"E8",
		x"B9" WHEN x"E9",
		x"F1" WHEN x"EA",
		x"09" WHEN x"EB",
		x"C5" WHEN x"EC",
		x"6E" WHEN x"ED",
		x"C6" WHEN x"EE",
		x"84" WHEN x"EF",
		x"18" WHEN x"F0",
		x"F0" WHEN x"F1",
		x"7D" WHEN x"F2",
		x"EC" WHEN x"F3",
		x"3A" WHEN x"F4",
		x"DC" WHEN x"F5",
		x"4D" WHEN x"F6",
		x"20" WHEN x"F7",
		x"79" WHEN x"F8",
		x"EE" WHEN x"F9",
		x"5F" WHEN x"FA",
		x"3E" WHEN x"FB",
		x"D7" WHEN x"FC",
		x"CB" WHEN x"FD",
		x"39" WHEN x"FE",
		x"48" WHEN x"FF",
		(OTHERS => '0') WHEN OTHERS;

END Behavioral;