LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ram IS
	PORT (
		CLK : IN STD_LOGIC;
		ROUNDKEY_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		WRITE_READ : IN STD_LOGIC;
		ROUNDKEY_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ram;

ARCHITECTURE Behavioral OF ram IS
	TYPE ram IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RAMDATA : ram;
BEGIN
	PROCESS (CLK) IS
	BEGIN
		IF (rising_edge(CLK)) THEN
			IF (WRITE_READ = '0') THEN
				-- Read operation
				ROUNDKEY_OUT <= RAMDATA(to_integer(unsigned(ADDRESS)));
			ELSE
				-- Write operation
				RAMDATA(to_integer(unsigned(ADDRESS))) <= ROUNDKEY_IN;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;