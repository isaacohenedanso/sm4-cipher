LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tribuffer IS
	PORT (
		INPT : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		EN : IN STD_LOGIC;
		OUTP : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END tribuffer;

ARCHITECTURE Behavioral OF tribuffer IS

BEGIN
	WITH EN SELECT
		OUTP <= INPT WHEN '1',
		"ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ" WHEN OTHERS;
END Behavioral;