LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SM4_TOP_MODEL_IMPLEMENTATION IS
    PORT (
        CLK, CLR, ENC_DEC : IN STD_LOGIC;
        MASTERKEY, INPUTTEXT : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
        OUTPUTTEXT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
    );
END SM4_TOP_MODEL_IMPLEMENTATION;

ARCHITECTURE BEHAVIORAL OF SM4_TOP_MODEL_IMPLEMENTATION IS
    COMPONENT Datapath IS
        PORT (
            INPUTTEXT, MASTERKEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
            OUTPUTTEXT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
            ENC_DEC, CLK, CLR, MKLOAD, ILOAD, XLOAD, MUXSEL1, MUXSEL2, MUXSEL3, MUXSEL4, WRITE_EN, OUTEN : IN STD_LOGIC;
            ILT32 : OUT STD_LOGIC
        );
    END COMPONENT;
    COMPONENT KeyExpansionCU IS
        PORT (
            CLR, CLK : IN STD_LOGIC;
            Ilt32 : IN STD_LOGIC;
            RST, WRITE_EN, MKLOAD, ILOAD, MUXSEL1, MUXSEL2, ROLLOVER : OUT STD_LOGIC
        );
    END COMPONENT;
    COMPONENT EncryptionDecryptionCU IS
        PORT (
            CLR, CLK : IN STD_LOGIC;
            ILT32 : IN STD_LOGIC;
            RST, WRITE_EN, XLOAD, ILOAD, MUXSEL3, OUTEN : OUT STD_LOGIC
        );
    END COMPONENT;
    COMPONENT mux3 IS
        PORT (
            INPT_A, INPT_B : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            SEL : IN STD_LOGIC;
            OUTP : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
        );
    END COMPONENT;

    SIGNAL IL32, MUX1, MUX2, SMUX3, ILD_KEY, ILD_ENC, W_KEY, W_ENC, ROLL, S_ROLL, MKLD, XLD, EN, RST_KEY, RST_ENC : STD_LOGIC;
    SIGNAL CTRL_KEY, CTRL_ENC, FROMMUX3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN

    S_ROLL <= NOT ROLL;
    CTRL_KEY <= RST_KEY & W_KEY & ILD_KEY;
    CTRL_ENC <= RST_ENC & W_ENC & ILD_ENC;

    Datapath0 : Datapath PORT MAP(
        INPUTTEXT => INPUTTEXT,
        MASTERKEY => MASTERKEY,
        OUTPUTTEXT => OUTPUTTEXT,
        ENC_DEC => ENC_DEC,
        CLK => CLK,
        CLR => FROMMUX3(2),
        MKLOAD => MKLD,
        ILOAD => FROMMUX3(0),
        XLOAD => XLD,
        MUXSEL1 => MUX1,
        MUXSEL2 => MUX2,
        MUXSEL3 => SMUX3,
        MUXSEL4 => ROLL,
        WRITE_EN => FROMMUX3(1),
        OUTEN => EN,
        ILT32 => IL32
    );
    KeyExpansionCU0 : KeyExpansionCU PORT MAP(
        CLR => CLR,
        CLK => CLK,
        RST => RST_KEY,
        ILT32 => IL32,
        WRITE_EN => W_KEY,
        MKLOAD => MKLD,
        ILOAD => ILD_KEY,
        MUXSEL1 => MUX1,
        MUXSEL2 => MUX2,
        ROLLOVER => ROLL
    );
    EncryptionDecryptionCU0 : EncryptionDecryptionCU PORT MAP(
        CLR => S_ROLL,
        CLK => CLK,
        RST => RST_ENC,
        ILT32 => IL32,
        WRITE_EN => W_ENC,
        XLOAD => XLD,
        ILOAD => ILD_ENC,
        MUXSEL3 => SMUX3,
        OUTEN => EN
    );
    mux3_0 : mux3 PORT MAP(
        INPT_A => CTRL_KEY,
        INPT_B => CTRL_ENC,
        SEL => ROLL,
        OUTP => FROMMUX3
    );
END BEHAVIORAL;