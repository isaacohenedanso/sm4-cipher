LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
-- 1 for enc 0 for dec
ENTITY CounterWithRam IS
	PORT (
		WRITE_EN, ENC_DEC, CLK, RST, ILOAD, MUXSEL4 : IN STD_LOGIC;
		ILT32 : OUT STD_LOGIC;
		ROUNDKEY_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ROUNDKEY_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		COUNT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END CounterWithRam;

ARCHITECTURE Behavioral OF CounterWithRam IS
	COMPONENT FF IS
		PORT (
			D, LOAD, CLK : IN STD_LOGIC;
			Q : OUT STD_LOGIC
		);
	END COMPONENT;
	COMPONENT mux1 IS
		PORT (
			SEL : IN STD_LOGIC;
			INPT_A, INPT_B : IN STD_LOGIC;
			OUTP : OUT STD_LOGIC
		);
	END COMPONENT;
	COMPONENT mux5 IS
		PORT (
			SEL : IN STD_LOGIC;
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT adder IS
		PORT (
			INPT : IN unsigned(5 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT substractor IS
		PORT (
			INPT : IN unsigned(4 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT ram IS
		PORT (
			CLK : IN STD_LOGIC;
			ROUNDKEY_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WRITE_READ : IN STD_LOGIC;
			ROUNDKEY_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT comparator_Ilt32 IS
		PORT (
			INPT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			OUTP : OUT STD_LOGIC
		);
	END COMPONENT;
	COMPONENT regi IS
		PORT (
			CLK, LOAD, RST : IN STD_LOGIC;
			D : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			Q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL FROMFF, FROMMUXAFTERFF : STD_LOGIC;
	SIGNAL FROMADDER, FROMREGI: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL FROMSUBTRACTOR, FROMMUX5_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN
	COUNT <= FROMREGI(4 DOWNTO 0);
	ff_E : FF PORT MAP(
		D => ENC_DEC,
		Q => FROMFF,
		LOAD => ILOAD,
		CLK => CLK
	);
	muxafterff : mux1 PORT MAP(
		SEL => MUXSEL4,
		INPT_A => FROMFF,
		INPT_B => '1',
		OUTP => FROMMUXAFTERFF
	);
	regi0 : regi PORT MAP(
		RST => RST,
		CLK => CLK,
		LOAD => ILOAD,
		D => FROMADDER,
		Q => FROMREGI
	);
	compare : comparator_Ilt32 PORT MAP(
		INPT => FROMREGI,
		OUTP => ILT32
	);
	add : adder PORT MAP(
		INPT => unsigned(FROMREGI),
		OUTP => FROMADDER
	);
	sub : substractor PORT MAP(
		INPT => unsigned(FROMREGI(4 DOWNTO 0)),
		OUTP => FROMSUBTRACTOR
	);
	mux5_0 : mux5 PORT MAP(
		SEL => FROMMUXAFTERFF,
		INPT_A => FROMSUBTRACTOR,
		INPT_B => FROMREGI(4 DOWNTO 0),
		OUTP => FROMMUX5_0
	);
	ramRK : ram PORT MAP(
		CLK => CLK,
		ROUNDKEY_IN => ROUNDKEY_IN,
		WRITE_READ => WRITE_EN,
		ADDRESS => FROMMUX5_0,
		ROUNDKEY_OUT => ROUNDKEY_OUT
	);
END Behavioral;