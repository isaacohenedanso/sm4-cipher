LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FF IS
	PORT (
		D, LOAD, CLK : IN STD_LOGIC;
		Q : OUT STD_LOGIC
	);
END FF;

ARCHITECTURE Behavioral OF FF IS

BEGIN
	PROCESS (CLK) IS
	BEGIN
		IF (rising_edge(CLK)) THEN
			IF (LOAD = '1') THEN
				Q <= D;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;