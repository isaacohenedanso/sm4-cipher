LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EncryptionDecryptionUnit IS
	PORT (
		XLOAD, CLK, MUXSEL3, OUTEN : IN STD_LOGIC;
		INPUTTEXT : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		ROUNDKEY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUTPUTTEXT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END EncryptionDecryptionUnit;

ARCHITECTURE Behavioral OF EncryptionDecryptionUnit IS
	COMPONENT reg128 IS
		PORT (
			CLK, LOAD : IN STD_LOGIC;
			D : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			Q : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_four IS
		PORT (
			INPT_A, INPT_B, INPT_C, INPT_D : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT sbox IS
		PORT (
			INPT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_two IS
		PORT (
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT tribuffer IS
		PORT (
			INPT : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			EN : IN STD_LOGIC;
			OUTP : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT mux128 IS
		PORT (
			SEL : IN STD_LOGIC;
			INPT_A, INPT_B : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT xor_five IS
		PORT (
			INPT_A, INPT_B, INPT_C, INPT_D, INPT_E : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL FROMREGX, NEXTINPT, RESHUFFLED, FROMMUX128, FROMREGO : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL FROMSBOXES, FROMXOR5_0, FROMXOR2_0, TOSBOXES, CIRC_SHIFT2, CIRC_SHIFT10, CIRC_SHIFT18, CIRC_SHIFT24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL FROMSBOX0, FROMSBOX1, FROMSBOX2, FROMSBOX3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
	FROMSBOXES <= FROMSBOX0 & FROMSBOX1 & FROMSBOX2 & FROMSBOX3;
	CIRC_SHIFT2 <= FROMSBOXES(29 DOWNTO 0) & FROMSBOXES(31 DOWNTO 30);
	CIRC_SHIFT10 <= FROMSBOXES(21 DOWNTO 0) & FROMSBOXES(31 DOWNTO 22);
	CIRC_SHIFT18 <= FROMSBOXES(13 DOWNTO 0) & FROMSBOXES(31 DOWNTO 14);
	CIRC_SHIFT24 <= FROMSBOXES(7 DOWNTO 0) & FROMSBOXES(31 DOWNTO 8);
	NEXTINPT <= FROMREGX(95 DOWNTO 0) & FROMXOR2_0;
	RESHUFFLED <= (NEXTINPT(31 DOWNTO 0) & NEXTINPT(63 DOWNTO 32) & NEXTINPT(95 DOWNTO 64) & NEXTINPT(127 DOWNTO 96));

	mux0 : mux128 PORT MAP(
		INPT_A => INPUTTEXT,
		INPT_B => NEXTINPT,
		SEL => MUXSEL3,
		OUTP => FROMMUX128
	);
	regX : reg128 PORT MAP(
		CLK => CLK,
		LOAD => XLOAD,
		D => FROMMUX128,
		Q => FROMREGX
	);
	xor4_0 : xor_four PORT MAP(
		INPT_A => FROMREGX(95 DOWNTO 64),
		INPT_B => FROMREGX(63 DOWNTO 32),
		INPT_C => FROMREGX(31 DOWNTO 0),
		INPT_D => ROUNDKEY,
		OUTP => TOSBOXES
	);
	sbox0 : sbox PORT MAP(
		INPT => TOSBOXES(31 DOWNTO 24),
		OUTP => FROMSBOX0
	);
	sbox1 : sbox PORT MAP(
		INPT => TOSBOXES(23 DOWNTO 16),
		OUTP => FROMSBOX1
	);
	sbox2 : sbox PORT MAP(
		INPT => TOSBOXES(15 DOWNTO 8),
		OUTP => FROMSBOX2
	);
	sbox3 : sbox PORT MAP(
		INPT => TOSBOXES(7 DOWNTO 0),
		OUTP => FROMSBOX3
	);
	xor5_0 : xor_five PORT MAP(
		INPT_A => FROMSBOXES,
		INPT_B => CIRC_SHIFT2,
		INPT_C => CIRC_SHIFT10,
		INPT_D => CIRC_SHIFT18,
		INPT_E => CIRC_SHIFT24,
		OUTP => FROMXOR5_0
	);
	xor2_0 : xor_two PORT MAP(
		INPT_A => FROMREGX(127 DOWNTO 96),
		INPT_B => FROMXOR5_0,
		OUTP => FROMXOR2_0
	);
	regO: reg128 port map(
		CLK => CLK,
		LOAD => XLOAD,
		D => RESHUFFLED,
		Q => FROMREGO			
		);
	buffer1 : tribuffer PORT MAP(
		INPT => FROMREGO,
		EN => OUTEN,
		OUTP => OUTPUTTEXT
	);
END Behavioral;