LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY rom IS
	PORT (
		INPT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		OUTP : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END rom;

ARCHITECTURE Behavioral OF rom IS
BEGIN
	WITH INPT SELECT
		OUTP <=
		x"00070E15" WHEN "00000",
		x"1C232A31" WHEN "00001",
		x"383F464D" WHEN "00010",
		x"545B6269" WHEN "00011",
		x"70777E85" WHEN "00100",
		x"8C939AA1" WHEN "00101",
		x"A8AFB6BD" WHEN "00110",
		x"C4CBD2D9" WHEN "00111",
		x"E0E7EEF5" WHEN "01000",
		x"FC030A11" WHEN "01001",
		x"181F262D" WHEN "01010",
		x"343B4249" WHEN "01011",
		x"50575E65" WHEN "01100",
		x"6C737A81" WHEN "01101",
		x"888F969D" WHEN "01110",
		x"A4ABB2B9" WHEN "01111",
		x"C0C7CED5" WHEN "10000",
		x"DCE3EAF1" WHEN "10001",
		x"F8FF060D" WHEN "10010",
		x"141B2229" WHEN "10011",
		x"30373E45" WHEN "10100",
		x"4C535A61" WHEN "10101",
		x"686F767D" WHEN "10110",
		x"848B9299" WHEN "10111",
		x"A0A7AEB5" WHEN "11000",
		x"BCC3CAD1" WHEN "11001",
		x"D8DFE6ED" WHEN "11010",
		x"F4FB0209" WHEN "11011",
		x"10171E25" WHEN "11100",
		x"2C333A41" WHEN "11101",
		x"484F565D" WHEN "11110",
		x"646B7279" WHEN "11111",
		x"00000000" WHEN OTHERS;
END Behavioral;